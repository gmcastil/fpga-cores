// Set to 1 to enable an ILA for the VGA core
`define ILA_VGA_CORE_ENABLE         1
// Set to 1 to enable an ILA just for the pattern generator
`define ILA_VGA_PATTERN_ENABLE      1

