// Set to 1 to enable an ILA for the VGA core
`define ILA_VGA_CORE    1

