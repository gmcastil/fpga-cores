`define   GND   1'b0
`define   VCC   1'b1

